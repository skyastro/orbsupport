  -36500.0  1.08634703e+11   2.0077
  -36450.0 1.103644407e+11   1.9938
  -36400.0 1.105242085e+11   1.9732
  -36350.0 1.088631027e+11   1.9764
  -36300.0 1.080415078e+11   1.9986
  -36250.0 1.094167024e+11   2.0017
  -36200.0 1.107321623e+11   1.9809
  -36150.0 1.099017839e+11   1.9666
  -36100.0 1.082340324e+11   1.9792
  -36050.0 1.084426127e+11   1.9957
  -36000.0 1.101819975e+11   1.9861
  -35950.0 1.106392361e+11   1.9639
  -35900.0 1.090956244e+11   1.9593
  -35850.0 1.080123083e+11   1.9765
  -35800.0 1.091745119e+11   1.9819
  -35750.0 1.106688527e+11   1.9629
  -35700.0 1.101160943e+11   1.9448
  -35650.0 1.083855013e+11   1.9506
  -35600.0   1.0828015e+11   1.9653
  -35550.0 1.099745851e+11   1.9576
  -35500.0 1.107157782e+11   1.9346
  -35450.0 1.093366698e+11   1.9253
  -35400.0 1.080270571e+11   1.9381
  -35350.0  1.08938346e+11   1.9432
  -35300.0 1.105661937e+11   1.9244
  -35250.0 1.103074113e+11   1.9038
  -35200.0 1.085684792e+11   1.9056
  -35150.0 1.081526824e+11   1.9182
  -35100.0 1.097484463e+11   1.9097
  -35050.0 1.107516048e+11   1.8849
  -35000.0 1.095786361e+11   1.8728
  -34950.0 1.080852577e+11   1.8837
  -34900.0 1.087157187e+11   1.8878
  -34850.0 1.104271858e+11   1.8663
  -34800.0 1.104700184e+11   1.8425
  -34750.0 1.087769587e+11   1.8428
  -34700.0 1.080644545e+11   1.8557
  -34650.0 1.095104684e+11   1.8453
  -34600.0 1.107456753e+11   1.8158
  -34550.0 1.098139908e+11   1.8004
  -34500.0 1.081849553e+11   1.8121
  -34450.0 1.085138017e+11   1.8174
  -34400.0 1.102559191e+11   1.7919
  -34350.0 1.105991031e+11   1.7619
  -34300.0  1.09004167e+11   1.7604
  -34250.0 1.080184217e+11   1.7767
  -34200.0 1.092679908e+11   1.7666
  -34150.0 1.106981617e+11   1.7302
  -34100.0 1.100355013e+11   1.7085
  -34050.0 1.083228151e+11   1.7215
  -34000.0 1.083391752e+11   1.7318
  -33950.0 1.100574751e+11   1.7036
  -33900.0 1.106908752e+11   1.6644
  -33850.0   1.0924281e+11   1.6583
  -33800.0 1.080161313e+11   1.6797
  -33750.0 1.090285903e+11   1.6740
  -33700.0  1.10610445e+11   1.6311
  -33650.0 1.102364447e+11   1.5993
  -33600.0  1.08494256e+11   1.6111
  -33550.0 1.081975882e+11   1.6294
  -33500.0 1.098378015e+11   1.6028
  -33450.0 1.107426562e+11   1.5537
  -33400.0 1.094853225e+11   1.5384
  -33350.0 1.080576605e+11   1.5631
  -33300.0 1.087998457e+11   1.5661
  -33250.0 1.104850841e+11   1.5206
  -33200.0 1.104107917e+11   1.4768
  -33150.0  1.08693628e+11   1.4825
  -33100.0 1.080937423e+11   1.5083
  -33050.0 1.096035572e+11   1.4884
  -33000.0 1.107529409e+11   1.4324
  -32950.0 1.097241166e+11   1.4048
  -32900.0 1.081416129e+11   1.4281
  -32850.0 1.085890911e+11   1.4411
  -32800.0  1.10325757e+11   1.3984
  -32750.0 1.105533642e+11   1.3440
  -32700.0 1.089144268e+11   1.3392
  -32650.0 1.080311088e+11   1.3689
  -32600.0  1.09361931e+11   1.3591
  -32550.0 1.107214308e+11   1.3011
  -32500.0 1.099518174e+11   1.2607
  -32450.0  1.08265175e+11   1.2773
  -32400.0  1.08403165e+11   1.2987
  -32350.0 1.101371748e+11   1.2636
  -32300.0 1.106599641e+11   1.2027
  -32250.0 1.091495306e+11   1.1849
  -32200.0 1.080117909e+11   1.2133
  -32150.0 1.091204347e+11   1.2138
  -32100.0 1.106490407e+11   1.1593
  -32050.0 1.101614815e+11   1.1090
  -32000.0 1.084242294e+11   1.1150
  -31950.0 1.082481654e+11   1.1402
  -31900.0 1.099249665e+11   1.1147
  -31850.0 1.107274736e+11   1.0528
  -31800.0 1.093914492e+11   1.0232
  -31750.0 1.080364387e+11   1.0451
  -31700.0  1.08886675e+11   1.0532
  -31650.0  1.10537879e+11   1.0059
  -31600.0 1.103467908e+11   0.9504
  -31550.0 1.086135163e+11   0.9445
  -31500.0 1.081292234e+11   0.9683
  -31450.0 1.096955359e+11   0.9521
  -31400.0 1.107539277e+11   0.8940
  -31350.0 1.096325747e+11   0.8558
  -31300.0 1.081042228e+11   0.8680
  -31250.0 1.086681107e+11   0.8792
  -31200.0 1.103911991e+11   0.8406
  -31150.0 1.105022207e+11   0.7850
  -31100.0 1.088268352e+11   0.7690
  -31050.0 1.080503054e+11   0.7869
  -31000.0 1.094558896e+11   0.7766
  -30950.0 1.107385583e+11   0.7250
  -30900.0 1.098654228e+11   0.6835
  -30850.0 1.082128681e+11   0.6860
  -30800.0 1.084718017e+11   0.6954
  -30750.0 1.102133241e+11   0.6636
  -30700.0 1.106231801e+11   0.6117
  -30650.0 1.090572741e+11   0.5900
  -30600.0 1.080140577e+11   0.6003
  -30550.0 1.092134405e+11   0.5914
  -30500.0 1.106818115e+11   0.5460
  -30450.0 1.100828586e+11   0.5054
  -30400.0 1.083587453e+11   0.5012
  -30350.0 1.083041609e+11   0.5060
  -30300.0 1.100095431e+11   0.4775
  -30250.0 1.107061231e+11   0.4304
  -30200.0 1.092974556e+11   0.4071
  -30150.0 1.080216994e+11   0.4113
  -30100.0 1.089757867e+11   0.4006
  -30050.0 1.105853376e+11   0.3588
  -30000.0 1.102783003e+11   0.3210
  -29950.0 1.085370151e+11   0.3141
  -29900.0  1.08170719e+11   0.3147
  -29850.0 1.097859787e+11   0.2860
  -29800.0 1.107486312e+11   0.2416
  -29750.0 1.095397881e+11   0.2194
  -29700.0 1.080729732e+11   0.2215
  -29650.0 1.087504738e+11   0.2088
  -29600.0 1.104519541e+11   0.1671
  -29550.0 1.104458981e+11   0.1303
  -29500.0 1.087418152e+11   0.1238
  -29450.0 1.080759145e+11   0.1240
  -29400.0 1.095494261e+11   0.0951
  -29350.0 1.107494696e+11   0.0497
  -29300.0 1.097767116e+11   0.0269
  -29250.0  1.08166156e+11   0.0302
  -29200.0 1.085447458e+11   0.0252
  -29150.0 1.102855806e+11   0.0321
  -29100.0 1.105806847e+11   0.0640
  -29050.0 1.089664805e+11   0.0700
  -29000.0 1.080229203e+11   0.0693
  -28950.0 1.093071659e+11   0.1002
  -28900.0 1.107086138e+11   0.1451
  -28850.0 1.100009304e+11   0.1682
  -28800.0 1.082981286e+11   0.1644
  -28750.0 1.083652953e+11   0.1743
  -28700.0 1.100911465e+11   0.2171
  -28650.0 1.106786978e+11   0.2572
  -28600.0 1.092037841e+11   0.2659
  -28550.0 1.080135172e+11   0.2609
  -28500.0 1.090667518e+11   0.2861
  -28450.0 1.106272508e+11   0.3338
  -28400.0  1.10205626e+11   0.3624
  -28350.0    1.084645e+11   0.3598
  -28300.0 1.082180208e+11   0.3630
  -28250.0  1.09874469e+11   0.4017
  -28200.0 1.107370746e+11   0.4460
  -28150.0 1.094461877e+11   0.4605
  -28100.0 1.080480216e+11   0.4539
  -28050.0  1.08835779e+11   0.4709
  -28000.0 1.105077523e+11   0.5168
  -27950.0 1.103846457e+11   0.5513
  -27900.0 1.086597794e+11   0.5537
  -27850.0 1.081078068e+11   0.5515
  -27800.0 1.096421038e+11   0.5822
  -27750.0 1.107541171e+11   0.6276
  -27700.0 1.096860905e+11   0.6497
  -27650.0  1.08125273e+11   0.6454
  -27600.0  1.08621638e+11   0.6536
  -27550.0 1.103536207e+11   0.6932
  -27500.0 1.105326643e+11   0.7322
  -27450.0  1.08877585e+11   0.7426
  -27400.0 1.080383338e+11   0.7384
  -27350.0 1.094011675e+11   0.7584
  -27300.0 1.107293305e+11   0.8005
  -27250.0 1.099160681e+11   0.8301
  -27200.0 1.082426808e+11   0.8324
  -27150.0 1.084312644e+11   0.8339
  -27100.0 1.101694072e+11   0.8632
  -27050.0 1.106453178e+11   0.9027
  -27000.0 1.091108779e+11   0.9224
  -26950.0 1.080119335e+11   0.9211
  -26900.0 1.091591345e+11   0.9311
  -26850.0 1.106634346e+11   0.9652
  -26800.0 1.101290935e+11   0.9989
  -26750.0 1.083963283e+11   1.0103
  -26700.0 1.082708917e+11   1.0100
  -26650.0 1.099606015e+11   1.0278
  -26600.0 1.107193082e+11   1.0627
  -26550.0 1.093522105e+11   1.0896
  -26500.0 1.080294941e+11   1.0955
  -26450.0 1.089236125e+11   1.0990
  -26400.0 1.105583471e+11   1.1221
  -26350.0 1.103187353e+11   1.1551
  -26300.0 1.085811278e+11   1.1756
  -26250.0 1.081458215e+11   1.1787
  -26200.0 1.097334928e+11   1.1868
  -26150.0 1.107524805e+11   1.2126
  -26100.0 1.095939772e+11   1.2425
  -26050.0 1.080904245e+11   1.2574
  -26000.0 1.087021009e+11   1.2600
  -25950.0 1.104171409e+11   1.2721
  -25900.0 1.104793305e+11   1.2991
  -25850.0 1.087910157e+11   1.3252
  -25800.0 1.080602203e+11   1.3355
  -25750.0 1.094950033e+11   1.3388
  -25700.0 1.107438712e+11   1.3541
  -25650.0  1.09828658e+11   1.3813
  -25600.0 1.081926786e+11   1.4032
  -25550.0 1.085017412e+11   1.4097
  -25500.0 1.102439725e+11   1.4145
  -25450.0 1.106061291e+11   1.4327
  -25400.0 1.090191786e+11   1.4590
  -25350.0 1.080169564e+11   1.4763
  -25300.0 1.092524945e+11   1.4801
  -25250.0 1.106937303e+11   1.4871
  -25200.0  1.10049047e+11   1.5074
  -25150.0 1.083328375e+11   1.5319
  -25100.0 1.083290673e+11   1.5442
  -25050.0 1.100439831e+11   1.5466
  -25000.0 1.106954095e+11   1.5562
  -24950.0 1.092582974e+11   1.5780
  -24900.0 1.080174842e+11   1.5992
  -24850.0 1.090135503e+11   1.6068
  -24800.0 1.106035153e+11   1.6094
  -24750.0 1.102484604e+11   1.6220
  -24700.0 1.085062456e+11   1.6440
  -24650.0 1.081897674e+11   1.6605
  -24600.0 1.098231708e+11   1.6645
  -24550.0  1.10744567e+11   1.6688
  -24500.0 1.095007982e+11   1.6840
  -24450.0  1.08061786e+11   1.7044
  -24400.0 1.087857414e+11   1.7155
  -24350.0 1.104758587e+11   1.7177
  -24300.0 1.104209189e+11   1.7247
  -24250.0 1.087071917e+11   1.7415
  -24200.0 1.080884692e+11   1.7584
  -24150.0 1.095882341e+11   1.7647
  -24100.0 1.107521726e+11   1.7673
  -24050.0 1.097390996e+11   1.7769
  -24000.0 1.081483724e+11   1.7934
  -23950.0 1.085763778e+11   1.8055
  -23900.0 1.103145075e+11   1.8089
  -23850.0 1.105613037e+11   1.8132
  -23800.0 1.089291247e+11   1.8246
  -23750.0 1.080285603e+11   1.8387
  -23700.0  1.09346389e+11   1.8461
  -23650.0 1.107180056e+11   1.8489
  -23600.0 1.099658483e+11   1.8553
  -23550.0 1.082743427e+11   1.8669
  -23500.0 1.083922577e+11   1.8771
  -23450.0 1.101242355e+11   1.8811
  -23400.0  1.10665483e+11   1.8848
  -23350.0 1.091648915e+11   1.8929
  -23300.0 1.080120527e+11   1.9029
  -23250.0 1.091051603e+11   1.9085
  -23200.0 1.106430583e+11   1.9111
  -23150.0 1.101741351e+11   1.9167
  -23100.0 1.084355008e+11   1.9253
  -23050.0 1.082394238e+11   1.9317
  -23000.0 1.099107257e+11   1.9336
  -22950.0  1.10730411e+11   1.9370
  -22900.0 1.094069871e+11   1.9443
  -22850.0  1.08039502e+11   1.9514
  -22800.0 1.088721528e+11   1.9531
  -22750.0 1.105295139e+11   1.9535
  -22700.0 1.103576881e+11   1.9589
  -22650.0 1.086265205e+11   1.9669
  -22600.0  1.08122938e+11   1.9702
  -22550.0 1.096804259e+11   1.9677
  -22500.0 1.107541983e+11   1.9689
  -22450.0 1.096478044e+11   1.9766
  -22400.0 1.081099846e+11   1.9835
  -22350.0 1.086548071e+11   1.9814
  -22300.0 1.103806969e+11   1.9765
  -22250.0 1.105110386e+11   1.9801
  -22200.0 1.088411484e+11   1.9897
  -22150.0 1.080466867e+11   1.9930
  -22100.0 1.094403751e+11   1.9851
  -22050.0 1.107361542e+11   1.9803
  -22000.0 1.098798749e+11   1.9875
  -21950.0 1.082211354e+11   1.9975
  -21900.0 1.084601491e+11   1.9943
  -21850.0 1.102009958e+11   1.9820
  -21800.0 1.106296594e+11   1.9800
  -21750.0 1.090724354e+11   1.9912
  -21700.0 1.080132272e+11   1.9986
  -21650.0 1.091980046e+11   1.9872
  -21600.0 1.106768025e+11   1.9734
  -21550.0 1.100960932e+11   1.9764
  -21500.0 1.083692429e+11   1.9908
  -21450.0 1.082945422e+11   1.9912
  -21400.0 1.099957571e+11   1.9722
  -21350.0 1.107100743e+11   1.9604
  -21300.0 1.093129829e+11   1.9702
  -21250.0 1.080236851e+11   1.9844
  -21200.0 1.089609166e+11   1.9744
  -21150.0 1.105778697e+11   1.9507
  -21100.0 1.102899193e+11   1.9445
  -21050.0 1.085493961e+11   1.9612
  -21000.0  1.08163453e+11   1.9698
  -20950.0 1.097711516e+11   1.9484
  -20900.0 1.107499396e+11   1.9242
  -20850.0  1.09555194e+11   1.9271
  -20800.0 1.080777083e+11   1.9479
  -20750.0 1.087366448e+11   1.9450
  -20700.0 1.104422459e+11   1.9143
  -20650.0 1.104555557e+11   1.8949
  -20600.0 1.087556746e+11   1.9088
  -20550.0 1.080712438e+11   1.9271
  -20500.0 1.095340115e+11   1.9093
  -20450.0 1.107480971e+11   1.8741
  -20400.0 1.097915189e+11   1.8652
  -20350.0 1.081734816e+11   1.8883
  -20300.0 1.085324055e+11   1.8960
  -20250.0 1.102739186e+11   1.8639
  -20200.0 1.105880959e+11   1.8309
  -20150.0 1.089813698e+11   1.8363
  -20100.0 1.080210017e+11   1.8619
  -20050.0 1.092916416e+11   1.8527
  -20000.0 1.107046002e+11   1.8109
  -19950.0 1.100146862e+11   1.7876
  -19900.0 1.083078001e+11   1.8074
  -19850.0 1.083548474e+11   1.8256
  -19800.0 1.100778779e+11   1.7979
  -19750.0 1.106836457e+11   1.7541
  -19700.0 1.092192276e+11   1.7468
  -19650.0 1.080144152e+11   1.7748
  -19600.0 1.090516052e+11   1.7765
  -19550.0 1.106207129e+11   1.7338
  -19500.0 1.102179147e+11   1.6972
  -19450.0 1.084761969e+11   1.7083
  -19400.0 1.082098107e+11   1.7337
  -19350.0  1.09859993e+11   1.7142
  -19300.0 1.107394151e+11   1.6644
  -19250.0 1.094616981e+11   1.6436
  -19200.0 1.080517061e+11   1.6687
  -19150.0 1.088214918e+11   1.6800
  -19100.0 1.104988812e+11   1.6409
  -19050.0    1.103951e+11   1.5945
  -19000.0 1.086731175e+11   1.5944
  -18950.0 1.081021077e+11   1.6225
  -18900.0 1.096268611e+11   1.6119
  -18850.0 1.107537821e+11   1.5609
  -18800.0  1.09701185e+11   1.5286
  -18750.0 1.081316201e+11   1.5466
  -18700.0 1.086086706e+11   1.5641
  -18650.0 1.103426773e+11   1.5313
  -18600.0 1.105409749e+11   1.4798
  -18550.0 1.088921308e+11   1.4685
  -18500.0 1.080353368e+11   1.4943
  -18450.0 1.093856281e+11   1.4911
  -18400.0 1.107263299e+11   1.4425
  -18350.0 1.099302827e+11   1.4025
  -18300.0  1.08251478e+11   1.4118
  -18250.0 1.084200393e+11   1.4313
  -18200.0  1.10156716e+11   1.4045
  -18150.0 1.106512407e+11   1.3516
  -18100.0 1.091261643e+11   1.3317
  -18050.0 1.080117393e+11   1.3529
  -18000.0 1.091437838e+11   1.3540
  -17950.0 1.106578555e+11   1.3086
  -17900.0 1.101419966e+11   1.2644
  -17850.0 1.084072834e+11   1.2663
  -17800.0 1.082617784e+11   1.2851
  -17750.0 1.099465427e+11   1.2622
  -17700.0 1.107226706e+11   1.2096
  -17650.0 1.093677529e+11   1.1844
  -17600.0 1.080321092e+11   1.2009
  -17550.0 1.089089364e+11   1.2033
  -17500.0 1.105503522e+11   1.1600
  -17450.0 1.103299399e+11   1.1140
  -17400.0 1.085938795e+11   1.1113
  -17350.0 1.081391227e+11   1.1284
  -17300.0 1.097184925e+11   1.1068
  -17250.0 1.107531846e+11   1.0539
  -17200.0 1.096092891e+11   1.0260
  -17150.0 1.080957611e+11   1.0400
  -17100.0   1.0868857e+11   1.0427
  -17050.0 1.104069646e+11   0.9992
  -17000.0 1.104885038e+11   0.9508
  -16950.0 1.088051479e+11   0.9458
  -16900.0 1.080561601e+11   0.9633
  -16850.0 1.094795217e+11   0.9425
  -16800.0 1.107418967e+11   0.8871
  -16750.0 1.098432665e+11   0.8556
  -16700.0 1.082005577e+11   0.8694
  -16650.0 1.084897944e+11   0.8748
  -16600.0 1.102319157e+11   0.8304
  -16550.0  1.10613001e+11   0.7771
  -16500.0 1.090342352e+11   0.7693
  -16450.0 1.080156709e+11   0.7897
  -16400.0 1.092370128e+11   0.7718
  -16350.0 1.106891344e+11   0.7126
  -16300.0 1.100625065e+11   0.6751
  -16250.0 1.083429964e+11   0.6887
  -16200.0 1.083190965e+11   0.6998
  -16150.0 1.100304056e+11   0.6565
  -16100.0 1.106997791e+11   0.5964
  -16050.0 1.092737987e+11   0.5829
  -16000.0 1.080190169e+11   0.6070
  -15950.0  1.08998556e+11   0.5959
  -15900.0 1.105964318e+11   0.5346
  -15850.0 1.102603653e+11   0.4879
  -15800.0 1.085183482e+11   0.4982
  -15750.0 1.081821026e+11   0.5167
  -15700.0  1.09808482e+11   0.4794
  -15650.0  1.10746307e+11   0.4133
  -15600.0 1.095162565e+11   0.3898
  -15550.0 1.080660852e+11   0.4147
  -15500.0 1.087717129e+11   0.4138
  -15450.0 1.104664948e+11   0.3555
  -15400.0 1.104309144e+11   0.2986
  -15350.0 1.087208416e+11   0.3007
  -15300.0 1.080833662e+11   0.3252
  -15250.0 1.095728827e+11   0.2987
  -15200.0 1.107512326e+11   0.2308
  -15150.0 1.097540351e+11   0.1942
  -15100.0 1.081552938e+11   0.2155
  -15050.0 1.085637682e+11   0.2251
  -15000.0 1.103031393e+11   0.1762
  -14950.0 1.105690944e+11   0.1115
  -14900.0 1.089438793e+11   0.1003
  -14850.0 1.080261902e+11   0.1269
  -14800.0 1.093308495e+11   0.1143
  -14750.0 1.107144129e+11   0.0575
  -14700.0 1.099798032e+11   0.0083
  -14650.0 1.082836549e+11   0.0183
  -14600.0  1.08381479e+11   0.0297
  -14550.0 1.101112007e+11   0.0337
  -14500.0 1.106708407e+11   0.0804
  -14450.0 1.091802784e+11   0.0993
  -14400.0 1.080124952e+11   0.0776
  -14350.0 1.090899197e+11   0.0801
  -14300.0 1.106369173e+11   0.1395
  -14250.0 1.101866871e+11   0.1901
  -14200.0 1.084468949e+11   0.1915
  -14150.0 1.082308315e+11   0.1705
  -14100.0 1.098964159e+11   0.1971
  -14050.0 1.107331795e+11   0.2593
  -14000.0 1.094225198e+11   0.2934
  -13950.0 1.080427422e+11   0.2805
  -13900.0 1.088576948e+11   0.2728
  -13850.0 1.105210039e+11   0.3177
  -13800.0 1.103684614e+11   0.3738
  -13750.0 1.086396216e+11   0.3891
  -13700.0  1.08116818e+11   0.3717
  -13650.0 1.096652759e+11   0.3834
  -13600.0 1.107542971e+11   0.4371
  -13550.0 1.096629982e+11   0.4802
  -13500.0 1.081159135e+11   0.4799
  -13450.0 1.086415966e+11   0.4687
  -13400.0 1.103700679e+11   0.4983
  -13350.0  1.10519714e+11   0.5513
  -13300.0 1.088555301e+11   0.5784
  -13250.0 1.080432438e+11   0.5698
  -13200.0  1.09424851e+11   0.5721
  -13150.0 1.107335805e+11   0.6131
  -13100.0 1.098942618e+11   0.6584
  -13050.0 1.082295546e+11   0.6708
  -13000.0 1.084486159e+11   0.6624
  -12950.0 1.101885626e+11   0.6794
  -12900.0 1.106359818e+11   0.7242
  -12850.0 1.090876348e+11   0.7580
  -12800.0 1.080125772e+11   0.7600
  -12750.0 1.091825903e+11   0.7587
  -12700.0  1.10671631e+11   0.7873
  -12650.0 1.101092357e+11   0.8294
  -12600.0  1.08379872e+11   0.8510
  -12550.0 1.082850653e+11   0.8488
  -12500.0 1.099818915e+11   0.8582
  -12450.0 1.107138591e+11   0.8930
  -12400.0 1.093285171e+11   0.9280
  -12350.0 1.080258498e+11   0.9390
  -12300.0  1.08946099e+11   0.9391
  -12250.0 1.105702511e+11   0.9585
  -12200.0 1.103014225e+11   0.9942
  -12150.0 1.085618844e+11   1.0198
  -12100.0 1.081563468e+11   1.0242
  -12050.0  1.09756273e+11   1.0308
  -12000.0 1.107510767e+11   1.0574
  -11950.0 1.095705758e+11   1.0897
  -11900.0 1.080826149e+11   1.1057
  -11850.0  1.08722898e+11   1.1085
  -11800.0 1.104324034e+11   1.1230
  -11750.0 1.104650772e+11   1.1528
  -11700.0 1.087696136e+11   1.1787
  -11650.0 1.080667456e+11   1.1870
  -11600.0 1.095185755e+11   1.1926
  -11550.0 1.107465535e+11   1.2140
  -11500.0 1.098062721e+11   1.2433
  -11450.0 1.081809655e+11   1.2610
  -11400.0 1.085201748e+11   1.2652
  -11350.0 1.102621428e+11   1.2765
  -11300.0 1.105953552e+11   1.3026
  -11250.0 1.089963091e+11   1.3278
  -11200.0 1.080192625e+11   1.3372
  -11150.0 1.092761268e+11   1.3414
  -11100.0 1.107004208e+11   1.3596
  -11050.0   1.1002836e+11   1.3873
  -11000.0 1.083176116e+11   1.4052
  -10950.0 1.083445331e+11   1.4083
  -10900.0 1.100645195e+11   1.4167
  -10850.0 1.106884303e+11   1.4409
  -10800.0 1.092346901e+11   1.4663
  -10750.0 1.080154935e+11   1.4753
  -10700.0 1.090364993e+11   1.4762
  -10650.0 1.106140192e+11   1.4911
  -10600.0 1.102300963e+11   1.5188
  -10550.0 1.084880109e+11   1.5380
  -10500.0 1.082017539e+11   1.5389
  -10450.0 1.098454543e+11   1.5422
  -10400.0 1.107415855e+11   1.5642
  -10350.0 1.094771963e+11   1.5915
  -10300.0 1.080555656e+11   1.6015
  -10250.0 1.088072757e+11   1.5975
  -10200.0 1.104898689e+11   1.6070
  -10150.0 1.104054257e+11   1.6347
  -10100.0 1.086865463e+11   1.6572
  -10050.0 1.080965768e+11   1.6569
  -10000.0 1.096115851e+11   1.6531
   -9950.0 1.107532755e+11   1.6709
   -9900.0 1.097162367e+11   1.7009
   -9850.0 1.081381312e+11   1.7141
   -9800.0 1.085958026e+11   1.7057
   -9750.0 1.103316115e+11   1.7071
   -9700.0 1.105491392e+11   1.7330
   -9650.0 1.089067383e+11   1.7604
   -9600.0 1.080325172e+11   1.7617
   -9550.0 1.093700861e+11   1.7501
   -9500.0 1.107231608e+11   1.7603
   -9450.0 1.099444258e+11   1.7916
   -9400.0  1.08260423e+11   1.8110
   -9350.0 1.084089389e+11   1.8011
   -9300.0 1.101439253e+11   1.7923
   -9250.0 1.106570041e+11   1.8124
   -9200.0 1.091414818e+11   1.8442
   -9150.0 1.080117258e+11   1.8515
   -9100.0 1.091284619e+11   1.8344
   -9050.0 1.106521161e+11   1.8335
   -9000.0 1.101548021e+11   1.8620
   -8950.0 1.084183649e+11   1.8887
   -8900.0 1.082528115e+11   1.8823
   -8850.0 1.099324104e+11   1.8641
   -8800.0 1.107258649e+11   1.8737
   -8750.0 1.093832951e+11   1.9068
   -8700.0 1.080349022e+11   1.9230
   -8650.0 1.088943198e+11   1.9053
   -8600.0 1.105422099e+11   1.8919
   -8550.0 1.103410238e+11   1.9123
   -8500.0 1.086067325e+11   1.9445
   -8450.0 1.081325871e+11   1.9468
   -8400.0 1.097034473e+11   1.9229
   -8350.0  1.10753717e+11   1.9189
   -8300.0   1.0962457e+11   1.9474
   -8250.0 1.081012667e+11   1.9729
   -8200.0 1.086751277e+11   1.9610
   -8150.0 1.103966583e+11   1.9375
   -8100.0 1.104975372e+11   1.9446
   -8050.0 1.088193531e+11   1.9770
   -8000.0 1.080522743e+11   1.9905
   -7950.0 1.094640256e+11   1.9679
   -7900.0 1.107397518e+11   1.9503
   -7850.0 1.098578144e+11   1.9680
   -7800.0 1.082085914e+11   1.9988
   -7750.0  1.08477963e+11   1.9976
   -7700.0 1.102197502e+11   1.9698
   -7650.0  1.10619718e+11   1.9617
   -7600.0 1.090493349e+11   1.9876
   -7550.0 1.080145656e+11   2.0109
   -7500.0 1.092215477e+11   1.9956
   -7450.0 1.106843744e+11   1.9686
   -7400.0 1.100758782e+11   1.9715
   -7350.0 1.083532905e+11   2.0014
   -7300.0 1.083092641e+11   2.0121
   -7250.0 1.100167442e+11   1.9865
   -7200.0 1.107039834e+11   1.9653
   -7150.0 1.092893118e+11   1.9791
   -7100.0 1.080207292e+11   2.0071
   -7050.0 1.089836094e+11   2.0028
   -7000.0 1.105891954e+11   1.9724
   -6950.0 1.102721581e+11   1.9605
   -6900.0 1.085305624e+11   1.9830
   -6850.0  1.08174595e+11   2.0027
   -6800.0 1.097937371e+11   1.9845
   -6750.0 1.107478763e+11   1.9549
   -6700.0 1.095316956e+11   1.9545
   -6650.0 1.080705575e+11   1.9811
   -6600.0 1.087577621e+11   1.9874
   -6550.0 1.104569937e+11   1.9592
   -6500.0 1.104407769e+11   1.9354
   -6450.0 1.087345758e+11   1.9467
   -6400.0 1.080784339e+11   1.9706
   -6350.0 1.095575047e+11   1.9615
   -6300.0 1.107501212e+11   1.9288
   -6250.0 1.097689213e+11   1.9152
   -6200.0  1.08162376e+11   1.9354
   -6150.0  1.08551264e+11   1.9494
   -6100.0 1.102916536e+11   1.9267
   -6050.0 1.105767356e+11   1.8955
   -6000.0 1.089586888e+11   1.8947
   -5950.0 1.080239986e+11   1.9177
   -5900.0 1.093153145e+11   1.9168
   -5850.0 1.107106531e+11   1.8849
   -5800.0 1.099936806e+11   1.8615
   -5750.0 1.082931105e+11   1.8730
   -5700.0 1.083708302e+11   1.8903
   -5650.0  1.10098072e+11   1.8735
   -5600.0 1.106760365e+11   1.8392
   -5550.0 1.091956892e+11   1.8282
   -5500.0 1.080131181e+11   1.8470
   -5450.0 1.090747148e+11   1.8511
   -5400.0 1.106306186e+11   1.8219
   -5350.0  1.10199136e+11   1.7923
   -5300.0 1.084584101e+11   1.7955
   -5250.0 1.082223896e+11   1.8126
   -5200.0 1.098820389e+11   1.8002
   -5150.0 1.107357786e+11   1.7650
   -5100.0 1.094380452e+11   1.7469
   -5050.0 1.080461586e+11   1.7605
   -5000.0 1.088433031e+11   1.7667
   -4950.0 1.105123501e+11   1.7395
   -4900.0 1.103791094e+11   1.7064
   -4850.0 1.086528179e+11   1.7034
   -4800.0  1.08110864e+11   1.7188
   -4750.0 1.096500876e+11   1.7084
   -4700.0 1.107542241e+11   1.6722
   -4650.0 1.096781541e+11   1.6497
   -4600.0 1.081220087e+11   1.6598
   -4550.0 1.086284811e+11   1.6664
   -4500.0 1.103593134e+11   1.6390
   -4450.0 1.105282456e+11   1.6028
   -4400.0 1.088699782e+11   1.5963
   -4350.0 1.080399772e+11   1.6112
   -4300.0 1.094093193e+11   1.6010
   -4250.0 1.107308374e+11   1.5620
   -4200.0 1.099085819e+11   1.5355
   -4150.0 1.082381244e+11   1.5445
   -4100.0 1.084372035e+11   1.5525
   -4050.0 1.101760259e+11   1.5234
   -4000.0 1.106421465e+11   1.4824
   -3950.0 1.091028702e+11   1.4728
   -3900.0 1.080121076e+11   1.4895
   -3850.0 1.091671997e+11   1.4807
   -3800.0 1.106662976e+11   1.4372
   -3750.0 1.101222847e+11   1.4049
   -3700.0 1.083906314e+11   1.4134
   -3650.0 1.082757314e+11   1.4257
   -3600.0 1.099679481e+11   1.3958
   -3550.0 1.107174769e+11   1.3474
   -3500.0  1.09344056e+11   1.3328
   -3450.0 1.080281931e+11   1.3528
   -3400.0 1.089313361e+11   1.3489
   -3350.0 1.105624827e+11   1.3011
   -3300.0 1.103128085e+11   1.2598
   -3250.0 1.085744782e+11   1.2658
   -3200.0 1.081494012e+11   1.2850
   -3150.0 1.097413448e+11   1.2581
   -3100.0 1.107520424e+11   1.2021
   -3050.0 1.095859313e+11   1.1784
   -3000.0 1.080876923e+11   1.2001
   -2950.0 1.087092354e+11   1.2046
   -2900.0 1.104224279e+11   1.1564
   -2850.0 1.104744618e+11   1.1047
   -2800.0 1.087836306e+11   1.1039
   -2750.0 1.080624204e+11   1.1291
   -2700.0 1.095031199e+11   1.1099
   -2650.0 1.107448391e+11   1.0491
   -2600.0 1.098209694e+11   1.0138
   -2550.0 1.081886067e+11   1.0326
   -2500.0 1.085080552e+11   1.0466
   -2450.0 1.102502546e+11   1.0032
   -2400.0 1.106024617e+11   0.9427
   -2350.0 1.090112964e+11   0.9307
   -2300.0 1.080177028e+11   0.9584
   -2250.0 1.092606236e+11   0.9503
   -2200.0  1.10696076e+11   0.8899
   -2150.0 1.100419503e+11   0.8425
   -2100.0 1.083275617e+11   0.8531
   -2050.0 1.083343539e+11   0.8748
   -2000.0 1.100510731e+11   0.8411
   -1950.0 1.106930509e+11   0.7762
   -1900.0 1.092501694e+11   0.7507
   -1850.0 1.080167519e+11   0.7752
   -1800.0 1.090214361e+11   0.7781
   -1750.0 1.106071705e+11   0.7240
   -1700.0 1.102421695e+11   0.6677
   -1650.0 1.084999405e+11   0.6661
   -1600.0 1.081938515e+11   0.6906
   -1550.0 1.098308548e+11   0.6687
   -1500.0 1.107435857e+11   0.6054
   -1450.0 1.094926802e+11   0.5676
   -1400.0 1.080595997e+11   0.5835
   -1350.0 1.087931325e+11   0.5943
   -1300.0 1.104807165e+11   0.5507
   -1250.0 1.104156216e+11   0.4909
   -1200.0 1.087000641e+11   0.4753
   -1150.0 1.080912148e+11   0.4967
   -1100.0 1.095962777e+11   0.4862
   -1050.0 1.107525971e+11   0.4302
   -1000.0 1.097312439e+11   0.3840
    -950.0 1.081448055e+11   0.3871
    -900.0 1.085830356e+11   0.4007
    -850.0  1.10320425e+11   0.3694
    -800.0 1.105571563e+11   0.3124
    -750.0 1.089214056e+11   0.2847
    -700.0 1.080298753e+11   0.2973
    -650.0 1.093545436e+11   0.2944
    -600.0 1.107198236e+11   0.2493
    -550.0 1.099584957e+11   0.2009
    -500.0 1.082695143e+11   0.1907
    -450.0 1.083979648e+11   0.2012
    -400.0 1.101310367e+11   0.1801
    -350.0 1.106626073e+11   0.1315
    -300.0 1.091568283e+11   0.0967
    -250.0 1.080118928e+11   0.0973
    -200.0 1.091131706e+11   0.0966
    -150.0 1.106462171e+11   0.0637
    -100.0 1.101675084e+11   0.0265
     -50.0 1.084295714e+11   0.0094
       0.0  1.08243992e+11   0.0000
      50.0 1.099182065e+11   0.0173
     100.0 1.107288908e+11   0.0595
     150.0  1.09398835e+11   0.0929
     200.0 1.080378726e+11   0.1000
     250.0 1.088797646e+11   0.1034
     300.0 1.105339212e+11   0.1310
     350.0 1.103519857e+11   0.1706
     400.0 1.086196851e+11   0.1935
     450.0 1.081262153e+11   0.1983
     500.0 1.096883591e+11   0.2122
     550.0 1.107540777e+11   0.2457
     600.0 1.096398178e+11   0.2779
     650.0 1.081069405e+11   0.2922
     700.0 1.086617759e+11   0.3004
     750.0 1.103862233e+11   0.3238
     800.0 1.105064296e+11   0.3570
     850.0 1.088336297e+11   0.3806
     900.0 1.080485635e+11   0.3911
     950.0 1.094485168e+11   0.4063
    1000.0 1.107374368e+11   0.4349
    1050.0    1.098723e+11   0.4636
    1100.0 1.082167786e+11   0.4801
    1150.0 1.084662484e+11   0.4919
    1200.0 1.102074776e+11   0.5140
    1250.0 1.106262793e+11   0.5432
    1300.0 1.090644755e+11   0.5655
    1350.0 1.080136405e+11   0.5782
    1400.0 1.092061012e+11   0.5945
    1450.0  1.10679451e+11   0.6210
    1500.0 1.100891604e+11   0.6474
    1550.0 1.083637184e+11   0.6640
    1600.0 1.082995715e+11   0.6765
    1650.0 1.100030006e+11   0.6978
    1700.0 1.107080219e+11   0.7255
    1750.0 1.093048348e+11   0.7475
    1800.0 1.080226209e+11   0.7601
    1850.0 1.089687124e+11   0.7748
    1900.0 1.105818069e+11   0.7999
    1950.0 1.102838372e+11   0.8266
    2000.0 1.085428864e+11   0.8439
    2050.0 1.081672456e+11   0.8546
    2100.0 1.097789378e+11   0.8728
    2150.0 1.107492745e+11   0.9000
    2200.0 1.095471135e+11   0.9240
    2250.0 1.080752024e+11   0.9368
    2300.0 1.087438906e+11   0.9477
    2350.0 1.104473565e+11   0.9695
    2400.0 1.104505053e+11   0.9973
    2450.0 1.087483926e+11   1.0173
    2500.0 1.080736731e+11   1.0264
    2550.0 1.095421023e+11   1.0391
    2600.0 1.107488386e+11   1.0642
    2650.0 1.097837562e+11   1.0912
    2700.0 1.081696181e+11   1.1065
    2750.0 1.085388669e+11   1.1130
    2800.0 1.102800519e+11   1.1287
    2850.0 1.105842262e+11   1.1565
    2900.0 1.089735511e+11   1.1814
    2950.0  1.08021986e+11   1.1911
    3000.0  1.09299786e+11   1.1965
    3050.0 1.107067268e+11   1.2162
    3100.0 1.100074787e+11   1.2461
    3150.0  1.08302708e+11   1.2669
    3200.0 1.083603128e+11   1.2707
    3250.0 1.100848512e+11   1.2775
    3300.0 1.106810699e+11   1.3022
    3350.0  1.09211122e+11   1.3325
    3400.0 1.080139215e+11   1.3464
    3450.0 1.090595476e+11   1.3456
    3500.0 1.106241628e+11   1.3565
    3550.0 1.102114801e+11   1.3863
    3600.0 1.084700449e+11   1.4140
    3650.0 1.082140995e+11   1.4192
    3700.0 1.098675964e+11   1.4168
    3750.0 1.107382082e+11   1.4342
    3800.0 1.094535613e+11   1.4678
    3850.0  1.08049751e+11   1.4890
    3900.0 1.088289795e+11   1.4856
    3950.0 1.105035535e+11   1.4856
    4000.0 1.103896307e+11   1.5108
    4050.0 1.086661077e+11   1.5448
    4100.0 1.081050771e+11   1.5559
    4150.0 1.096348632e+11   1.5468
    4200.0 1.107539793e+11   1.5532
    4250.0 1.096932702e+11   1.5854
    4300.0 1.081282693e+11   1.6151
    4350.0 1.086154623e+11   1.6145
    4400.0 1.103484346e+11   1.6046
    4450.0 1.105366325e+11   1.6201
    4500.0 1.088844909e+11   1.6565
    4550.0 1.080368873e+11   1.6767
    4600.0  1.09393782e+11   1.6662
    4650.0 1.107279253e+11   1.6608
    4700.0 1.099228332e+11   1.6859
    4750.0 1.082468437e+11   1.7215
    4800.0 1.084259136e+11   1.7285
    4850.0 1.101633875e+11   1.7131
    4900.0 1.106481528e+11   1.7164
    4950.0 1.091181396e+11   1.7492
    5000.0 1.080118187e+11   1.7778
    5050.0 1.091518348e+11   1.7718
    5100.0 1.106608028e+11   1.7575
    5150.0 1.101352385e+11   1.7713
    5200.0 1.084015195e+11   1.8073
    5250.0  1.08266542e+11   1.8237
    5300.0 1.099539285e+11   1.8088
    5350.0 1.107209273e+11   1.8007
    5400.0 1.093595978e+11   1.8244
    5450.0 1.080307149e+11   1.8574
    5500.0 1.089166296e+11   1.8598
    5550.0 1.105545655e+11   1.8417
    5600.0 1.103240758e+11   1.8433
    5650.0  1.08587176e+11   1.8736
    5700.0 1.081426173e+11   1.8973
    5750.0 1.097263688e+11   1.8878
    5800.0 1.107528365e+11   1.8725
    5850.0 1.096012588e+11   1.8845
    5900.0 1.080929399e+11   1.9161
    5950.0 1.086956586e+11   1.9267
    6000.0 1.104123203e+11   1.9102
    6050.0  1.10483708e+11   1.9021
    6100.0 1.087977236e+11   1.9229
    6150.0 1.080582688e+11   1.9493
    6200.0 1.094876468e+11   1.9468
    6250.0  1.10742954e+11   1.9292
    6300.0 1.098356089e+11   1.9304
    6350.0 1.081964042e+11   1.9558
    6400.0 1.084960486e+11   1.9719
    6450.0 1.102382555e+11   1.9599
    6500.0 1.106094146e+11   1.9462
    6550.0 1.090263296e+11   1.9565
    6600.0 1.080163229e+11   1.9808
    6650.0  1.09245134e+11   1.9845
    6700.0 1.106915663e+11   1.9682
    6750.0 1.100554552e+11   1.9615
    6800.0 1.083376491e+11   1.9785
    6850.0 1.083243109e+11   1.9960
    6900.0 1.100375402e+11   1.9888
    6950.0  1.10697507e+11   1.9731
    7000.0 1.092656637e+11   1.9749
    7050.0 1.080181903e+11   1.9941
    7100.0 1.090064176e+11   2.0009
    7150.0 1.106001676e+11   1.9869
    7200.0 1.102541327e+11   1.9759
    7250.0  1.08511984e+11   1.9853
    7300.0 1.081861047e+11   2.0008
    7350.0 1.098161963e+11   1.9965
    7400.0 1.107454153e+11   1.9806
    7450.0 1.095081479e+11   1.9769
    7500.0 1.080638078e+11   1.9906
    7550.0  1.08779064e+11   1.9973
    7600.0 1.104714252e+11   1.9847
    7650.0 1.104256863e+11   1.9716
    7700.0 1.087136689e+11   1.9758
    7750.0 1.080860225e+11   1.9880
    7800.0 1.095809409e+11   1.9838
    7850.0 1.107517472e+11   1.9675
    7900.0 1.097462046e+11   1.9608
    7950.0 1.081516421e+11   1.9708
    8000.0 1.085703714e+11   1.9757
    8050.0 1.103091188e+11   1.9619
    8100.0 1.105650253e+11   1.9468
    8150.0 1.089361307e+11   1.9486
    8200.0 1.080274115e+11   1.9591
    8250.0 1.093390026e+11   1.9530
    8300.0 1.107163188e+11   1.9337
    8350.0 1.099724907e+11   1.9245
    8400.0 1.082787509e+11   1.9338
    8450.0 1.083871184e+11   1.9381
    8500.0 1.101180518e+11   1.9208
    8550.0 1.106680496e+11   1.9013
    8600.0 1.091722018e+11   1.9017
    8650.0 1.080122405e+11   1.9137
    8700.0  1.09097912e+11   1.9062
    8750.0 1.106401592e+11   1.8810
    8800.0 1.101801139e+11   1.8675
    8850.0 1.084409013e+11   1.8779
    8900.0 1.082353211e+11   1.8849
    8950.0 1.099039327e+11   1.8637
    9000.0  1.10731748e+11   1.8366
    9050.0 1.094143707e+11   1.8341
    9100.0 1.080410201e+11   1.8502
    9150.0 1.088652727e+11   1.8447
    9200.0 1.105254871e+11   1.8126
    9250.0 1.103628243e+11   1.7908
    9300.0 1.086327355e+11   1.8012
    9350.0 1.081200085e+11   1.8146
    9400.0 1.096732299e+11   1.7928
    9450.0 1.107542667e+11   1.7560
    9500.0 1.096550307e+11   1.7462
    9550.0 1.081127819e+11   1.7663
    9600.0 1.086485163e+11   1.7676
    9650.0 1.103756607e+11   1.7309
    9700.0 1.105151799e+11   1.6976
    9750.0 1.088479757e+11   1.7039
    9800.0 1.080450283e+11   1.7250
    9850.0 1.094329975e+11   1.7077
    9900.0  1.10734952e+11   1.6622
    9950.0 1.098867213e+11   1.6412
   10000.0 1.082251182e+11   1.6619
   10050.0 1.084546523e+11   1.6728
   10100.0 1.101950992e+11   1.6364
   10150.0 1.106326841e+11   1.5913
   10200.0 1.090796552e+11   1.5887
   10250.0 1.080128958e+11   1.6153
   10300.0 1.091906753e+11   1.6069
   10350.0 1.106743647e+11   1.5569
   10400.0 1.101023515e+11   1.5227
   10450.0 1.083742787e+11   1.5386
   10500.0   1.0829002e+11   1.5588
   10550.0 1.099891765e+11   1.5281
   10600.0 1.107118941e+11   1.4744
   10650.0 1.093203657e+11   1.4592
   10700.0 1.080246917e+11   1.4864
   10750.0  1.08953867e+11   1.4885
   10800.0 1.105742673e+11   1.4397
   10850.0 1.102954014e+11   1.3938
   10900.0 1.085553186e+11   1.4001
   10950.0 1.081600554e+11   1.4259
   11000.0  1.09764086e+11   1.4043
   11050.0 1.107505014e+11   1.3469
   11100.0 1.095625082e+11   1.3188
   11150.0 1.080800191e+11   1.3413
   11200.0 1.087301005e+11   1.3524
   11250.0 1.104375844e+11   1.3092
   11300.0 1.104600983e+11   1.2555
   11350.0   1.0876229e+11   1.2500
   11400.0 1.080690843e+11   1.2764
   11450.0 1.095266773e+11   1.2645
   11500.0 1.107473847e+11   1.2085
   11550.0  1.09798538e+11   1.1700
   11600.0 1.081770191e+11   1.1836
   11650.0 1.085265784e+11   1.1997
   11700.0 1.102683356e+11   1.1646
   11750.0 1.105915653e+11   1.1084
   11800.0 1.089884645e+11   1.0916
   11850.0 1.080201527e+11   1.1136
   11900.0  1.09284266e+11   1.1089
   11950.0 1.107026344e+11   1.0581
   12000.0 1.100211958e+11   1.0139
   12050.0 1.083124462e+11   1.0174
   12100.0 1.083499282e+11   1.0334
   12150.0 1.100715397e+11   1.0058
   12200.0 1.106859403e+11   0.9514
   12250.0 1.092265748e+11   0.9267
   12300.0 1.080149053e+11   0.9413
   12350.0 1.090444201e+11   0.9400
   12400.0 1.106175508e+11   0.8954
   12450.0 1.102237181e+11   0.8498
   12500.0 1.084817976e+11   0.8448
   12550.0  1.08205962e+11   0.8572
   12600.0 1.098530904e+11   0.8343
   12650.0 1.107404679e+11   0.7840
   12700.0 1.094690662e+11   0.7556
   12750.0 1.080535187e+11   0.7630
   12800.0 1.088147259e+11   0.7609
   12850.0 1.104946151e+11   0.7208
   12900.0  1.10400024e+11   0.6771
   12950.0 1.086794891e+11   0.6677
   13000.0 1.080994578e+11   0.6750
   13050.0 1.096196044e+11   0.6530
   13100.0 1.107535627e+11   0.6060
   13150.0 1.097083446e+11   0.5778
   13200.0 1.081346944e+11   0.5811
   13250.0 1.086025419e+11   0.5762
   13300.0 1.103374328e+11   0.5373
   13350.0 1.105448737e+11   0.4954
   13400.0 1.088990663e+11   0.4851
   13450.0 1.080339745e+11   0.4897
   13500.0 1.093782411e+11   0.4664
   13550.0 1.107248446e+11   0.4200
   13600.0  1.09937014e+11   0.3923
   13650.0 1.082557113e+11   0.3949
   13700.0 1.084147476e+11   0.3890
   13750.0 1.101506488e+11   0.3490
   13800.0     1.10654e+11   0.3065
   13850.0 1.091334411e+11   0.2963
   13900.0 1.080117103e+11   0.3016
   13950.0 1.091364975e+11   0.2782
   14000.0 1.106551474e+11   0.2296
   14050.0 1.101480954e+11   0.2003
   14100.0 1.084125348e+11   0.2040
   14150.0 1.082574981e+11   0.2007
   14200.0 1.099398346e+11   0.1604
   14250.0 1.107242098e+11   0.1138
   14300.0 1.093751403e+11   0.1019
   14350.0 1.080334146e+11   0.1101
   14400.0 1.089019815e+11   0.0919
   14450.0 1.105465004e+11   0.0429
   14500.0 1.103352233e+11   0.0054
   14550.0 1.085999761e+11   0.0084
   14600.0 1.081359959e+11   0.0175
   14650.0 1.097113469e+11   0.0389
   14700.0 1.107534591e+11   0.0799
   14750.0 1.096165562e+11   0.0955
   14800.0 1.080983569e+11   0.0856
   14850.0 1.086821696e+11   0.1022
   14900.0 1.104020821e+11   0.1516
   14950.0  1.10492815e+11   0.1893
   15000.0 1.088118907e+11   0.1904
   15050.0 1.080542913e+11   0.1842
   15100.0  1.09472158e+11   0.2173
   15150.0 1.107408984e+11   0.2681
   15200.0 1.098501888e+11   0.2918
   15250.0 1.082043569e+11   0.2833
   15300.0 1.084841564e+11   0.2896
   15350.0 1.102261469e+11   0.3351
   15400.0  1.10616213e+11   0.3793
   15450.0 1.090414069e+11   0.3880
   15500.0 1.080151231e+11   0.3788
   15550.0 1.092296599e+11   0.4012
   15600.0 1.106868924e+11   0.4511
   15650.0 1.100688732e+11   0.4832
   15700.0 1.083478724e+11   0.4806
   15750.0 1.083144057e+11   0.4794
   15800.0 1.100239226e+11   0.5154
   15850.0 1.107017981e+11   0.5620
   15900.0 1.092811708e+11   0.5803
   15950.0 1.080198083e+11   0.5732
   16000.0 1.089914457e+11   0.5849
   16050.0 1.105930113e+11   0.6282
   16100.0 1.102659846e+11   0.6662
   16150.0 1.085241399e+11   0.6730
   16200.0 1.081785145e+11   0.6686
   16250.0 1.098014806e+11   0.6927
   16300.0 1.107470742e+11   0.7367
   16350.0 1.095235973e+11   0.7641
   16400.0 1.080681894e+11   0.7637
   16450.0 1.087650722e+11   0.7670
   16500.0  1.10461996e+11   0.7996
   16550.0 1.104356187e+11   0.8395
   16600.0 1.087273591e+11   0.8568
   16650.0 1.080810005e+11   0.8545
   16700.0 1.095655766e+11   0.8670
   16750.0 1.107507257e+11   0.9033
   16800.0 1.097611168e+11   0.9365
   16850.0   1.0815864e+11   0.9460
   16900.0 1.085578117e+11   0.9462
   16950.0 1.102976946e+11   0.9664
   17000.0  1.10572745e+11   1.0024
   17050.0 1.089509116e+11   1.0282
   17100.0 1.080251262e+11   1.0329
   17150.0  1.09323465e+11   1.0380
   17200.0 1.107126467e+11   1.0632
   17250.0  1.09986409e+11   1.0966
   17300.0 1.082881314e+11   1.1156
   17350.0 1.083764012e+11   1.1185
   17400.0 1.101049722e+11   1.1286
   17450.0 1.106733305e+11   1.1562
   17500.0 1.091876003e+11   1.1859
   17550.0 1.080127688e+11   1.1993
   17600.0 1.090826881e+11   1.2023
   17650.0 1.106339431e+11   1.2167
   17700.0 1.101926171e+11   1.2451
   17750.0 1.084523531e+11   1.2705
   17800.0 1.082268002e+11   1.2794
   17850.0 1.098895907e+11   1.2840
   17900.0  1.10734436e+11   1.3019
   17950.0 1.094299001e+11   1.3299
   18000.0 1.080443441e+11   1.3503
   18050.0  1.08850846e+11   1.3560
   18100.0 1.105169086e+11   1.3631
   18150.0 1.103735382e+11   1.3838
   18200.0 1.086458821e+11   1.4100
   18250.0 1.081139673e+11   1.4250
   18300.0 1.096580615e+11   1.4291
   18350.0 1.107542838e+11   1.4394
   18400.0 1.096702067e+11   1.4620
   18450.0 1.081187899e+11   1.4849
   18500.0 1.086353508e+11   1.4948
   18550.0 1.103649718e+11   1.4990
   18600.0 1.105237871e+11   1.5128
   18650.0 1.088623892e+11   1.5358
   18700.0 1.080416691e+11   1.5539
   18750.0 1.094174695e+11   1.5598
   18800.0 1.107322978e+11   1.5660
   18850.0 1.099010767e+11   1.5828
   18900.0 1.082336091e+11   1.6042
   18950.0 1.084431764e+11   1.6166
   19000.0 1.101826166e+11   1.6208
   19050.0 1.106389316e+11   1.6302
   19100.0 1.090948719e+11   1.6487
   19150.0 1.080123315e+11   1.6661
   19200.0  1.09175272e+11   1.6735
   19250.0 1.106691161e+11   1.6785
   19300.0 1.101154498e+11   1.6914
   19350.0 1.083849699e+11   1.7091
   19400.0 1.082806109e+11   1.7210
   19450.0 1.099752737e+11   1.7255
   19500.0 1.107155995e+11   1.7335
   19550.0 1.093359023e+11   1.7485
   19600.0 1.080269413e+11   1.7629
   19650.0 1.089390752e+11   1.7693
   19700.0 1.105665774e+11   1.7739
   19750.0  1.10306849e+11   1.7853
   19800.0 1.085678572e+11   1.8002
   19850.0 1.081530254e+11   1.8092
   19900.0 1.097491836e+11   1.8121
   19950.0 1.107515571e+11   1.8194
   20000.0 1.095778777e+11   1.8332
   20050.0  1.08085007e+11   1.8449
   20100.0 1.087163935e+11   1.8481
   20150.0 1.104276785e+11   1.8508
   20200.0 1.104695549e+11   1.8618
   20250.0 1.087762664e+11   1.8759
   20300.0 1.080646682e+11   1.8818
   20350.0 1.095112317e+11   1.8808
   20400.0 1.107457599e+11   1.8863
   20450.0 1.098132649e+11   1.9006
   20500.0 1.081845779e+11   1.9117
   20550.0 1.085144003e+11   1.9108
   20600.0 1.102565062e+11   1.9088
   20650.0 1.105987521e+11   1.9188
   20700.0 1.090034268e+11   1.9344
   20750.0 1.080184987e+11   1.9394
   20800.0 1.092687565e+11   1.9327
   20850.0 1.106983763e+11   1.9333
   20900.0 1.100348301e+11   1.9481
   20950.0 1.083223237e+11   1.9616
   21000.0  1.08339678e+11   1.9583
   21050.0 1.100581392e+11   1.9492
   21100.0 1.106906469e+11   1.9551
   21150.0 1.092420455e+11   1.9729
   21200.0 1.080160692e+11   1.9806
   21250.0 1.090293342e+11   1.9693
   21300.0 1.106107833e+11   1.9618
   21350.0 1.102358484e+11   1.9740
   21400.0 1.084936668e+11   1.9920
   21450.0 1.081979785e+11   1.9904
   21500.0 1.098385226e+11   1.9737
   21550.0 1.107425575e+11   1.9714
   21600.0 1.094845578e+11   1.9895
   21650.0 1.080574613e+11   2.0034
   21700.0 1.088005442e+11   1.9912
   21750.0 1.104855361e+11   1.9734
   21800.0 1.104102881e+11   1.9785
   21850.0 1.086929604e+11   2.0003
   21900.0 1.080940071e+11   2.0054
   21950.0 1.096043132e+11   1.9840
   22000.0 1.107529744e+11   1.9697
   22050.0 1.097233754e+11   1.9834
   22100.0 1.081412832e+11   2.0045
   22150.0 1.085897216e+11   1.9973
   22200.0 1.103263095e+11   1.9707
   22250.0 1.105529682e+11   1.9639
   22300.0 1.089137024e+11   1.9851
   22350.0 1.080312393e+11   1.9999
   22400.0 1.093626987e+11   1.9797
   22450.0 1.107215956e+11   1.9531
   22500.0 1.099511225e+11   1.9565
   22550.0  1.08264726e+11   1.9821
   22600.0  1.08403707e+11   1.9847
   22650.0 1.101378113e+11   1.9542
   22700.0 1.106596873e+11   1.9331
   22750.0 1.091487726e+11   1.9478
   22800.0 1.080117826e+11   1.9715
   22850.0 1.091211899e+11   1.9585
   22900.0 1.106493321e+11   1.9230
   22950.0  1.10160854e+11   1.9121
   23000.0 1.084236759e+11   1.9365
   23050.0  1.08248601e+11   1.9506
   23100.0 1.099256681e+11   1.9225
   23150.0 1.107273241e+11   1.8885
   23200.0 1.093906817e+11   1.8914
   23250.0  1.08036292e+11   1.9197
   23300.0 1.088873939e+11   1.9176
   23350.0 1.105382884e+11   1.8788
   23400.0 1.103462494e+11   1.8532
   23450.0 1.086128766e+11   1.8705
   23500.0  1.08129538e+11   1.8936
   23550.0 1.096962811e+11   1.8729
   23600.0 1.107539099e+11   1.8305
   23650.0 1.096318216e+11   1.8193
   23700.0 1.081039426e+11   1.8464
   23750.0 1.086687701e+11   1.8553
   23800.0 1.103917145e+11   1.8186
   23850.0 1.105017815e+11   1.7811
   23900.0 1.088261301e+11   1.7871
   23950.0 1.080504887e+11   1.8149
   24000.0 1.094566556e+11   1.8038
   24050.0 1.107386726e+11   1.7582
   24100.0 1.098647074e+11   1.7335
   24150.0 1.082124637e+11   1.7544
   24200.0 1.084723803e+11   1.7716
   24250.0 1.102139302e+11   1.7409
   24300.0 1.106228561e+11   1.6957
   24350.0 1.090565263e+11   1.6894
   24400.0 1.080141034e+11   1.7166
   24450.0 1.092142034e+11   1.7145
   24500.0 1.106820546e+11   1.6700
   24550.0 1.100822026e+11   1.6351
   24600.0 1.083582303e+11   1.6472
   24650.0 1.083046396e+11   1.6684
   24700.0 1.100102219e+11   1.6444
   24750.0 1.107059236e+11   1.5959
   24800.0 1.092966889e+11   1.5790
   24850.0 1.080216059e+11   1.6022
   24900.0 1.089765225e+11   1.6062
   24950.0 1.105857025e+11   1.5648
   25000.0 1.102777235e+11   1.5235
   25050.0 1.085364065e+11   1.5268
   25100.0  1.08171082e+11   1.5483
   25150.0 1.097867096e+11   1.5299
   25200.0 1.107485622e+11   1.4809
   25250.0 1.095390266e+11   1.4565
   25300.0 1.080727438e+11   1.4741
   25350.0 1.087511589e+11   1.4809
   25400.0   1.1045243e+11   1.4427
   25450.0 1.104454177e+11   1.3982
   25500.0 1.087411328e+11   1.3947
   25550.0 1.080761496e+11   1.4144
   25600.0 1.095501868e+11   1.3989
   25650.0 1.107495329e+11   1.3500
   25700.0 1.097759789e+11   1.3211
   25750.0 1.081657984e+11   1.3346
   25800.0 1.085453581e+11   1.3422
   25850.0 1.102861536e+11   1.3050
   25900.0 1.105803147e+11   1.2580
   25950.0 1.089657464e+11   1.2507
   26000.0 1.080230197e+11   1.2695
   26050.0 1.093079328e+11   1.2551
   26100.0 1.107088077e+11   1.2045
   26150.0 1.100002489e+11   1.1721
   26200.0 1.082976546e+11   1.1839
   26250.0 1.083658147e+11   1.1928
   26300.0 1.100917995e+11   1.1550
   26350.0 1.106784492e+11   1.1043
   26400.0 1.092030219e+11   1.0940
   26450.0 1.080134775e+11   1.1141
   26500.0 1.090675009e+11   1.1013
   26550.0 1.106275696e+11   1.0473
   26600.0 1.102050164e+11   1.0100
   26650.0 1.084639254e+11   1.0212
   26700.0 1.082184303e+11   1.0341
   26750.0 1.098751823e+11   0.9961
   26800.0 1.107369546e+11   0.9392
   26850.0 1.094454213e+11   0.9244
   26900.0 1.080478442e+11   0.9475
   26950.0 1.088364864e+11   0.9398
   27000.0 1.105081868e+11   0.8824
   27050.0 1.103841261e+11   0.8369
   27100.0 1.086591231e+11   0.8459
   27150.0 1.081080926e+11   0.8655
   27200.0 1.096428558e+11   0.8311
   27250.0 1.107541291e+11   0.7672
   27300.0 1.096853439e+11   0.7440
   27350.0 1.081249638e+11   0.7690
   27400.0  1.08622281e+11   0.7698
   27450.0  1.10354158e+11   0.7126
   27500.0 1.105322501e+11   0.6573
   27550.0 1.088768682e+11   0.6601
   27600.0 1.080384864e+11   0.6861
   27650.0 1.094019349e+11   0.6598
   27700.0 1.107294743e+11   0.5916
   27750.0 1.099153643e+11   0.5570
   27800.0 1.082422501e+11   0.5799
   27850.0  1.08431822e+11   0.5908
   27900.0 1.101700314e+11   0.5391
   27950.0 1.106450211e+11   0.4748
   28000.0 1.091101237e+11   0.4668
   28050.0 1.080119478e+11   0.4960
   28100.0 1.091598934e+11   0.4817
   28150.0 1.106637059e+11   0.4146
   28200.0 1.101284537e+11   0.3674
   28250.0 1.083957906e+11   0.3826
   28300.0 1.082713456e+11   0.4021
   28350.0 1.099612939e+11   0.3615
   28400.0 1.107191378e+11   0.2928
   28450.0 1.093514429e+11   0.2705
   28500.0 1.080293695e+11   0.2976
   28550.0 1.089243388e+11   0.2956
   28600.0 1.105587381e+11   0.2363
   28650.0 1.103181788e+11   0.1789
   28700.0 1.085805007e+11   0.1818
   28750.0 1.081461565e+11   0.2054
   28800.0 1.097342324e+11   0.1788
   28850.0 1.107524412e+11   0.1135
   28900.0 1.095932202e+11   0.0754
   28950.0 1.080901653e+11   0.0952
   29000.0 1.087027715e+11   0.1025
   29050.0 1.104176401e+11   0.0615
   29100.0 1.104788739e+11   0.0225
   29150.0 1.087903197e+11   0.0201
   29200.0 1.080604254e+11   0.0074
   29250.0 1.094957675e+11   0.0239
   29300.0 1.107439643e+11   0.0785
   29350.0 1.098279349e+11   0.1161
   29400.0 1.081922935e+11   0.1097
   29450.0 1.085023342e+11   0.0968
   29500.0 1.102445651e+11   0.1354
   29550.0 1.106057857e+11   0.1924
   29600.0 1.090184362e+11   0.2148
   29650.0 1.080170245e+11   0.2008
   29700.0 1.092532595e+11   0.2060
   29750.0 1.106939531e+11   0.2556
   29800.0   1.1004838e+11   0.3019
   29850.0 1.083323393e+11   0.3084
   29900.0 1.083295633e+11   0.2974
   29950.0 1.100446515e+11   0.3211
   30000.0 1.106951894e+11   0.3724
   30050.0 1.092575322e+11   0.4040
   30100.0 1.080174131e+11   0.4008
   30150.0  1.09014292e+11   0.4012
   30200.0 1.106038612e+11   0.4375
   30250.0 1.102478695e+11   0.4826
   30300.0 1.085056507e+11   0.5002
   30350.0   1.0819015e+11   0.4957
   30400.0 1.098238948e+11   0.5101
   30450.0 1.107444766e+11   0.5510
   30500.0 1.095000342e+11   0.5857
   30550.0 1.080615782e+11   0.5933
   30600.0 1.087864363e+11   0.5949
   30650.0 1.104763175e+11   0.6204
   30700.0 1.104204218e+11   0.6592
   30750.0 1.087065198e+11   0.6829
   30800.0 1.080887257e+11   0.6867
   30850.0 1.095889916e+11   0.6974
   30900.0 1.107522145e+11   0.7286
   30950.0 1.097383607e+11   0.7612
   31000.0 1.081480348e+11   0.7761
   31050.0 1.085770033e+11   0.7816
   31100.0 1.103150659e+11   0.8008
   31150.0  1.10560915e+11   0.8326
   31200.0 1.089283974e+11   0.8576
   31250.0  1.08028682e+11   0.8675
   31300.0 1.093471566e+11   0.8782
   31350.0 1.107181787e+11   0.9028
   31400.0 1.099651571e+11   0.9314
   31450.0 1.082738865e+11   0.9493
   31500.0 1.083927934e+11   0.9584
   31550.0 1.101248768e+11   0.9749
   31600.0 1.106652142e+11   1.0013
   31650.0 1.091641322e+11   1.0248
   31700.0 1.080120356e+11   1.0377
   31750.0 1.091059139e+11   1.0490
   31800.0 1.106433575e+11   1.0700
   31850.0 1.101735125e+11   1.0954
   31900.0 1.084349412e+11   1.1135
   31950.0 1.082398521e+11   1.1238
   32000.0 1.099114307e+11   1.1386
   32050.0 1.107302699e+11   1.1621
   32100.0 1.094062198e+11   1.1847
   32150.0 1.080393466e+11   1.1978
   32200.0 1.088728685e+11   1.2078
   32250.0 1.105299305e+11   1.2262
   32300.0 1.103571528e+11   1.2505
   32350.0 1.086258759e+11   1.2690
   32400.0 1.081232446e+11   1.2781
   32450.0 1.096811731e+11   1.2897
   32500.0  1.10754189e+11   1.3115
   32550.0 1.096470531e+11   1.3347
   32600.0 1.081096961e+11   1.3480
   32650.0 1.086554619e+11   1.3547
   32700.0 1.103812186e+11   1.3695
   32750.0 1.105106065e+11   1.3937
   32800.0 1.088404399e+11   1.4139
   32850.0 1.080468613e+11   1.4215
   32900.0 1.094411416e+11   1.4280
   32950.0 1.107362769e+11   1.4470
   33000.0 1.098791626e+11   1.4721
   33050.0 1.082207235e+11   1.4871
   33100.0 1.084607219e+11   1.4899
   33150.0 1.102016071e+11   1.4987
   33200.0 1.106293431e+11   1.5220
   33250.0 1.090716857e+11   1.5458
   33300.0  1.08013264e+11   1.5538
   33350.0 1.091987665e+11   1.5537
   33400.0 1.106770537e+11   1.5670
   33450.0 1.100954417e+11   1.5937
   33500.0 1.083687213e+11   1.6133
   33550.0  1.08295014e+11   1.6137
   33600.0 1.099964399e+11   1.6140
   33650.0 1.107098831e+11   1.6334
   33700.0 1.093122159e+11   1.6614
   33750.0 1.080235828e+11   1.6733
   33800.0 1.089616498e+11   1.6675
   33850.0 1.105782421e+11   1.6719
   33900.0 1.102893482e+11   1.6975
   33950.0 1.085487821e+11   1.7231
   34000.0 1.081638082e+11   1.7250
   34050.0 1.097718851e+11   1.7165
   34100.0  1.10749879e+11   1.7281
   34150.0 1.095544337e+11   1.7583
   34200.0 1.080774704e+11   1.7770
   34250.0 1.087373258e+11   1.7691
   34300.0 1.104427286e+11   1.7626
   34350.0 1.104550819e+11   1.7826
   34400.0 1.087549882e+11   1.8137
   34450.0 1.080714705e+11   1.8218
   34500.0 1.095347734e+11   1.8070
   34550.0 1.107481689e+11   1.8069
   34600.0 1.097907888e+11   1.8345
   34650.0 1.081731161e+11   1.8617
   34700.0 1.085330124e+11   1.8573
   34750.0 1.102744973e+11   1.8407
   34800.0 1.105877334e+11   1.8498
   34850.0 1.089806333e+11   1.8825
   34900.0 1.080210923e+11   1.9003
   34950.0 1.092924081e+11   1.8849
   35000.0 1.107048023e+11   1.8719
   35050.0 1.100140087e+11   1.8911
   35100.0 1.083073191e+11   1.9241
   35150.0 1.083553603e+11   1.9287
   35200.0 1.100785353e+11   1.9065
   35250.0 1.106834052e+11   1.9015
   35300.0 1.092184644e+11   1.9296
   35350.0 1.080143666e+11   1.9570
   35400.0 1.090523523e+11   1.9474
   35450.0 1.106210395e+11   1.9243
   35500.0 1.102173102e+11   1.9301
   35550.0 1.084756164e+11   1.9634
   35600.0 1.082102126e+11   1.9794
   35650.0 1.098607094e+11   1.9583
   35700.0 1.107393035e+11   1.9399
   35750.0 1.094609324e+11   1.9570
   35800.0   1.0805152e+11   1.9899
   35850.0 1.088221958e+11   1.9909
   35900.0 1.104993226e+11   1.9636
   35950.0 1.103945867e+11   1.9543
   36000.0 1.086724566e+11   1.9810
   36050.0 1.081023853e+11   2.0066
   36100.0 1.096276148e+11   1.9927
   36150.0 1.107538027e+11   1.9652
   36200.0 1.097004405e+11   1.9677
   36250.0 1.081313027e+11   1.9998
   36300.0 1.086093087e+11   2.0121
   36350.0 1.103432206e+11   1.9867
   36400.0 1.105405679e+11   1.9647
   36450.0  1.08891411e+11   1.9798
   36500.0 1.080354807e+11   2.0104
